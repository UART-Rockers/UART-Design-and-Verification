

class uart_config_class;
static virtual uart_intf svif;
static mailbox gen2bfm =new();
static mailbox mon2sbd =new();
static mailbox mon2sbd1 =new();
static string Operated_mode;
static string testname;

endclass
 
